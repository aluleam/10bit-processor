    Mac OS X            	   2  �     �                                    ATTR���  �  H   �                 H     com.apple.quarantine   _     com.apple.TextEncoding     n     com.apple.provenance   y     com.apple.lastuseddate#PS 4   �   y  7com.apple.metadata:kMDLabel_kvvvmagl5khnneff2fecvox3ey   0086;67448a43;TextEdit;utf-8;134217984  �<�B�T�@�Dg    ��]
    ��I���_^������Fܾ�n�g�OA΍�+�+ܲ�n�p0S1�_XC�L��g��8ˤ,�f�>���ы� 
�SÜ?���O��|�j�gu� �O�\0 �����B�[�.���YQ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             This resource fork intentionally left blank                                                                                                                                                                                                                            ��