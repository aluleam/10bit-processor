    Mac OS X            	   2  �     �                                    ATTR���_  �  H   �                 H     com.apple.quarantine   _     com.apple.TextEncoding     n     com.apple.provenance   y     com.apple.lastuseddate#PS 4   �   y  7com.apple.metadata:kMDLabel_kvvvmagl5khnneff2fecvox3ey   0086;67448a11;TextEdit;utf-8;134217984  �<�B�T��Dg    �"    ���Y�_X�.]�/p�~� S�*&�v�0e�9x&��T�K���'_O�@�t8�`�1�!�S�D�B�pc�Dc���J!�gո��_	�/_��5�ʘ������'n�D��A䭔��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             This resource fork intentionally left blank                                                                                                                                                                                                                            ��