    Mac OS X            	   2  �     �                                    ATTR���8  �  H   �                 H     com.apple.quarantine   _     com.apple.TextEncoding     n     com.apple.provenance   y     com.apple.lastuseddate#PS 4   �   y  7com.apple.metadata:kMDLabel_kvvvmagl5khnneff2fecvox3ey   0086;67448a35;TextEdit;utf-8;134217984  �<�B�T�3�Dg    �D�-    򺄭�(�T����[VM�ٔ��4���_�UW#�Y�J�6�����^d��Ӆ��f4��D��|Pe吔��:0@�!o������������P��*�����8�O{($��i%+���sE�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             This resource fork intentionally left blank                                                                                                                                                                                                                            ��